library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library lib_VHDL;
use lib_VHDL.present_library.all;


entity key_Schedule is
   port(
	reset		: in std_logic;
	clk		: in std_logic;

	key  		: in std_logic_vector(79 downto 0);       	
        round_Counter	: in std_logic_vector(4 downto 0);
	CNT		: in CNT_key_Schedule;

	round_Key	: out std_logic_vector(63 downto 0)
	);
	
end key_Schedule;

architecture A of key_Schedule is

	component register_80_bits is
   		port(	reg_in  	: in  std_logic_vector(79 downto 0);
			enable		: in  std_logic;
			reset		: in  std_logic;
			clk		: in  std_logic;
			reg_out		: out std_logic_vector(79 downto 0));
	end component;

	component s_Box_4_Bits is
  		port( 	s_Box_In  	: in  std_logic_vector(3 downto 0);
        		s_Box_Out	: out std_logic_vector(3 downto 0));
	end component;

signal s_Box_Out : std_logic_vector(3 downto 0);
signal add_Round_Counter_Out : std_logic_vector(4 downto 0);
signal mux_Out : std_logic_vector(79 downto 0);
signal register_Out : std_logic_vector(79 downto 0);
signal register_Rotation : std_logic_vector(79 downto 0);

begin

	REG: register_80_bits port map (mux_Out, CNT.write, reset, clk, register_Out);

	SBOX: s_Box_4_Bits port map (register_Rotation(79 downto 76), s_Box_Out);

	ADD: add_Round_Counter_Out <= register_Rotation(19 downto 15) XOR round_Counter;

	ROT: register_Rotation(79 downto 0) <= register_Out(18 downto 0) & register_Out(79 downto 19);

	round_Key <= register_Out(79 downto 16);

	process (CNT.mux, clk, s_Box_Out, add_Round_Counter_Out, register_Rotation)
	begin
		if (CNT.mux = '1') then
			mux_Out <= key;
		else
			mux_Out <= s_Box_Out & register_Rotation(75 downto 20) & add_Round_Counter_Out & register_Rotation(14 downto 0);
		end if;
	end process;
			
	

end A;

































