library IEEE;
use IEEE.STD_LOGIC_1164.all;
library lib_VHDL;


package present_library is

	constant ROUND_KEY_SIZE : natural := 64;
	constant ROUND_COUNTER_SIZE : natural := 5;

	type CNT_key_Schedule is
	record
		mux 		: STD_LOGIC;
		write 		: STD_LOGIC;
	end record;

	type CNT_block_Cypher is
	record
		text_In 		: STD_LOGIC;
		write 		: STD_LOGIC;
		text_Out	: STD_LOGIC;
	end record;

	type CNT_memory is
	record
		write 		: STD_LOGIC;
	end record;

	type CNT is
	record
		memory 		: CNT_memory;
		key_Schedule 	: CNT_key_Schedule;
		block_Cypher 	: CNT_block_Cypher;
	end record;

	type MODE_TYPE is (CRYP, DECRYP);

	type KEY_SIZE is (K_80, K_128);



end present_library ;
