work.register_WIDTH_bits(A) :64:
work.s_Box_4_Bits(A) rtlc_no_parameters
